

module if_fifo_read(
);
endmodule
